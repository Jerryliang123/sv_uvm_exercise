interface ahb_inter;
  bit hclk=0;
  bit hreset=0;  
  bit[1:0] htrans;
endinterface  