/* properties: 
   methods:
    1.  
    2.
    3.
*/
class ReceiverBase;
    
    function new();
        ;
        
    endfunction

endclass //ReceiverBase

/* properties: 
   methods:
    1. 
    2.
    3.
*/
class Receiver;
    function new();
        
    endfunction //new()
endclass //Receiver